BZh91AY&SY�^Y� 
�_�Pyc��g߰����`
�=���   �dP���(I�P�35@��@����i���$��M@4a0�@���� L� �h0  bh�A&��D���@��   @���a2dɑ��4�# C �$�4�mL�O)�jd4�4 i�M5�
�@���̞��dI^У�	�����?�$��s�!��L`g���:���ڬ%)kE�-T���R �Qeݨ]Z� �H�Ԉ�"r�E�D�ԈQh��
`*����-z�Rf�]a���:h��Ģ��$C"��fّ�C+�'�uHY��5KJ�q9nX��1�ŉ��.�A$��V��"TқAcw#)B�N�51��M��VVܛ�V��\ˌf�gsYf)�
���>�����l�Ā�YtnnQ�IF�rn�Ō�T�@^B�` �W;�H���Ƙ��.|w)a�L�U�m�Σ7Nú����nȸ�n��̼ܻ�Swl��;��cwn!��n�̫�ښ�Ǘ�����׻;��ѧ�v63s72�nw^�R%IrdL�a19dK� ���B�2�C��ׄ4��KPBX�p))��HQT�W�Q�Kf3D�vxD3�$QE�6+�{��s��ÀvYH\/.sY��W����65p��3��E�\�
F�FF,m]r�89���p��u���2���,4�i�.=>�Ab��	�l� Zk�*��i���p
��g���M�zy� $�zn�\KP�j�́}���M09g�zy�%c��u �|X�:�<�H���ΐs�T)�K�;9�yE�,0�6�!�G��c[�x���g����5�]w�˱�:���{�*z�z�u $��؂�0�+!�s�R�D��s��j��pN�3�D��b�����M����Υ�o��Ƃ�2�b�
4A9ճ�ɑ��e
�x3���=#m鎤3G��������Ka���9!�챤3G�*�d+�����f�q�O�Ǟ`L0�I6ڒ�����q�(�求�2����6r���`�/]t����yޕy�F���ʍ�	u=;�gD�+g:�؉A&�l0�0��s|#lc��j���ʆ���yQ��^��nCcs��S��B�ah��!i�1D���^��0���a�������$��2m��t�>Fł,&\Aes�.�@Rx�6�k��������ې�����J�@���m�[L��@�E��a�ٜ�#zj0Ma�`Aڧaɭ��uɗ��KBFTڪ�
�&��OG�>Q��@����G;�3�;~�k�ʕ������Y�[Ɉ>F��C�J�u�K.�D�͜��[;ОN�5�w�%�I�㽎=�:���PQ����E��f���x��wݸx0n1r4�^9�c�E~�=��xA �}�I2Q��v��7����>��Q-rű�1b^RA��i``X�b��$0c0"@�`�����i!A
���,0 ��,0�J�IRI�`�*	E��%�,4�2!c1CDǬ�7�`�����.�`{k�l�?Y�W��3w�3�1ܕ��5Kob�v�ȧ�-B)n��s�pbV��C�P����?Gpwr{m����A@}�HP�M/o9������[�����!����L���d�i{���20`1l�?��HFeDF�3�/Y	��3�%�zs��L��h3zt��P��S���u�>a ��b��G�>8���x�!�˕�٘��47-�}��k
F⃶���Xx���ު	u��:	%8dmq�AJ	!C��9��d�&ާL����f�~AK����y��u�ù6]2x���� �Yx��\����n�tD`�C����,����2��yX)�3���I
�z1-Q,qw�.���|8<��8�=〼ZJ��&��.�c�H�1�AY%q'�v��>��vt�F  �@�u�0:��@�;G�ǔK�I�q�4i\I:������99�;�m��C�ɛHtk/�ĵ��-�����h�D9�n�5�
Csq��f8��n`�Q`rͣ^������;/$�R$�
�I�EVSAJ>e�`B�r���5�/�]��BCUyf�