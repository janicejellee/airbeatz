BZh91AY&SY��w a߀Pyc��g߰����`�n=��Zh(QB�7�<� &����yM�T �h��dO
��F�#��h4�j���*A� �0���  ��UL�4�Ѡb��4�d`LM&L�LM2100E!5<@��cR�&��C5  z��S~r	�1���$k���$dE��0�j3�8�"�Y�?�v�&h�%K:b��M���z�7�/ey�$-��@"У�TD����e�(R�N�kJ�n�dE�Il@�2��E��7FV�eE�e�V�F(Ֆ����������6 D���e$r��'E+u:-��ݕ:�-,����nX��e#�e����i����^ �=]A��V�U�_��Z���L]d���cbMp�6��sL�:�ˌ�2æ܍;w��N�Ƕ�����:�jj\ʇ�n�U&�s�
���)��I�y�4a�mɭ�5"��L�*eI�9�P��v��gaj���7-���TVɣ���*�.xX�0�C�l��G�3�����/��O�++~�ƎSF�tKo�&\�8�����䙙��V�U�l���.�����}u��r���
 L   �� p �H 
��jNs( �@ P`�
 A9ړ   �� 	 p�N��Ųd�ɓ��t��?�u8q�X>
���6I�Q�igҊ"';�e�e�g�e,����&�����m��m���s��v��C��?�ZJ��&tX��+C�"K�gM�n�b��1��{Ud�]h�X�wiź�����ԶY�Vw�j�0�uWV`J���!A(�  @(P�m���8���򗁭^ӳ}`E� DD/��#�lHҳ�T��r��]��U�|���?z��L;����y��߅�(�b�w�3Jț��{ƴ��jt�	f!Ly�fR};3BM��V�@�$��(S����oz<*�b�N����O����wfF1&�m$O�`�  P�(� $(B+����Lm|o���lo�x��q�x��o�W����    Uw�n:��e�7Nt*i�T�${a�6��
`Re����
��!?%OT���M���B�>HT�b�⩯�]Z�9��bbF�"ς�PX��V�uP���Ǝ̀��A$+?dF.��x�#mBP�5��P%?�$��@(�  I>� әW+����qN>���   ��;���v�vQ�Y1�/�K�1��H��A��b�4H@��H�K�,��:� �v��h�,QfW�AT[A�u1�z�eq5��L��)ex��(7v(���U��)ZB){���n��	$�JB(� �@	B��P:�/����Y�^/�^�ңcc��E   C�;�CXh\�s4��8�K}�G���)L�X_�O�����;L,$�Mj�P����t�^0�'z_m�&�\��IN-:��gd/��\�gB���V/!F��V]��-ͼ�9f��;�d|�et���5�&��)JWZԼ���� �  M��8�X���5����K`D,�S�I��˪�6{j�җDA���fd�G�T�H�(��s��F��]���T5G3զ�u1�ə���dAF������   ���9�^+��w�:Ьg�G	̺�����(M�ҍ��i�-ڌU�Vw�Y�/`�lF��හGh�+S������	B���M�����9�bCF7�cq�`7v��;�    ��0��{�g����ߏH��:HG��z�S�����˘���8���)�L��:��E�;�"�[
"�^���&/�u4+�Zɩºv�����m}g�9�   �[�95�reW�X�k�2�o/.;青1c�Ҧv�Q�[s��и�xg��s�V�����8�6t��MO+���p�|�jK�>֞��[vF=�(�L�c8�g�j��YbY�y   ,\ŭ�݆���v*�����R!r��}Q3�UۉWE�+��4�`�C�B�©�1�S���_ʻ4E���A��,�b��_KL�]lU�ue�sԾ^�2y�nB!�[m�d�#>~�3�ŒK�	�2�����\��c8R���,��𩱑�1k�d�3�#(\T��2�IqS�!�IK
QJ)E,�Y*B�����E,)dRR��AQK
TR�Y��J���ZZ(����)d=��f.�d��aM,�t^�`�$&N췝x$��?_�[mw�Z����mJ/�ٟ*��IB�Ut����.�Ɗ��I(gZ��¹��FWY������L�Dv��4���=�{�c�&�Rđ��0�#t�r�ܹ4���1���f؇��D{X��'���d�r�������VEL8��{�a�ɯfvI�i����'��?��͕��}�>�3�Ĉwʏ
���e�����Ň��tG�GA����Qe$Ya	q��~Z�Sh�Wso\[8kuL�	�/s�O�����Rđu:��\�����~.���ї��d��z5D�ws���:L��]���iմ�"68Z^G��ڹ�ӳ���n�vDH�">׸Xx�n�8�ms:f���82��~�K4p��dH�F��g��1#��14bYv1{���=Uڬk�L����g��GfF��~>}�/wS�$���f<��b���ۖ���v�V�!�,=]������',��>�tmg$��&�#����"8��6ƌ͑�登t��͒a]�����.7N���5,�����M�F���{N��Z�[wgDhσ���ta]m�x�Y�r��zzf����tg%���5n߾J��n�����f�^jВ[�jwm�6�g�y:e�YI4�k���.�p�!��.�