BZh91AY&SY숳� !_�Pxc��g߰����P�s�t .'"�Z�$I Bx%<���hz&&�i��@�@"��zF � i�� �	M=R$L�&�@bbh��@4i��&�&	��0`��$�dҞ�b��O)� �2�z�4�ytD�bBa!D-$�jυ�<@��x���ǅ�*������9ZSɶxuw�+w%���*��������vݭ⵷e����6z��m�$� ���L�Ah,��{�9���L�CAJ�D��ieⰤg�~�����n@��l��%m��ݹ�^ɛe4c|D�Y\�T������k���r]�"��j����NL���E��/UW.�v-O�{}G�  tA=}g�n���z�h�h�/煦��2���M�%1!�l*��("U���+�"��L� k���N�íA$����U�Y�EΡ�mš��T^��A�n&a)"L wb�m$A ��N�l[h�B�J����	9-��l79����EHa\�u�&�������F�^s@��(9"�#��+\gu"E�MrY��C�ˑoS���E���KY��lK*r�r�,��rI'���D�X����H)ۅ�>�4_���$�0..ET6'�9�[�Y,�i��k0�I��.f3�~���n[�S[�qn-�yn=nN���8�.�\���dd8v6랪x����m� xyv�XG7���`9U�$��u Bѡ
HHJ	p�P"(Ԩ76v�T��q�ar�km�S�k3�l��뎇G1U,�áH����ô�1$|i?�j�t�e���.���}ӫ���k�=�x�����N͟��w����X�3y��Â\jw�\�O��S�(�-��,gV{�+	!��Z�5o�*��S��MS4��'����۝M�(d��Wd�a&�5�I�H�MY���
�Ḱ����i��1��ñn�Ry
�Sn�����{��=�� qy%�v��Uؒ#m�-p�A��a�a|��\�S_��8�d�T��,���3V��e(�ƤC�W��JN��k�m�e:�mf�WF���T�eݾ}�$B��cG���j�K%��^ 9�l���fܤ�2@�`UΟÿ��ǘ��ղj����c*C۷/M
B��+2ݬz������Z�dj��\������u�p_�W]�-Q���j�H&8���Pˌ.�̪�Si�<��.��]����-���s���Z70:2i�n��D��h�It�~t>�gAӰ��Q�"�1�ߍ���=3|�8�[/��<��.�p�!�g8